library verilog;
use verilog.vl_types.all;
entity xor_32_bits_TB is
end xor_32_bits_TB;
