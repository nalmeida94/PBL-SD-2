library verilog;
use verilog.vl_types.all;
entity TB_shifter_right_32_bits is
end TB_shifter_right_32_bits;
