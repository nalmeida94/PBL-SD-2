library verilog;
use verilog.vl_types.all;
entity TB_or_32_bits is
end TB_or_32_bits;
