library verilog;
use verilog.vl_types.all;
entity TB_xor_32_bits is
end TB_xor_32_bits;
