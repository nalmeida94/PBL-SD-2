library verilog;
use verilog.vl_types.all;
entity TB_shifter_left_32_bits is
end TB_shifter_left_32_bits;
