library verilog;
use verilog.vl_types.all;
entity TB_subtrator_32_bits is
end TB_subtrator_32_bits;
