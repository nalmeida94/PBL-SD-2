library verilog;
use verilog.vl_types.all;
entity TB_and_32_bits is
end TB_and_32_bits;
