library verilog;
use verilog.vl_types.all;
entity TB_not_32_bits is
end TB_not_32_bits;
