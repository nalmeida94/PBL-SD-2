library verilog;
use verilog.vl_types.all;
entity TB_somador_32_bits is
end TB_somador_32_bits;
